module test(
  input        clock,
  input  [7:0] a,
  input  [7:0] b
);
endmodule
